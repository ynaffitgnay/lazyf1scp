module M0(__clk,__in_read,__in_vid,__in_data,__in_valid,__out_data,__out_valid);
	input wire __clk;
	input wire __in_read;
	input wire[13:0] __in_vid;
	input wire[63:0] __in_data;
	input wire __in_valid;
	output wire[63:0] __out_data;
	output wire __out_valid;
	(*shreg_extract = "no"*) reg[238:0] __read_buf[3:2];
	(*shreg_extract = "no"*) reg[238:0] __write_buf[3:2];
	(*shreg_extract = "no"*) reg[63:0] __in_buf[3:2];
	reg[63:0] __out_buf[1:0];
	reg[63:0] __out;
	(*shreg_extract = "no"*) reg __out_valid_buf[3:0];
	wire[238:0] __read;
	wire[238:0] __write;
	wire[63:0] __in;
	wire __wait;
	reg[63:0] __var[238:0];
	reg __feof[63:0];
	(*non_volatile*) reg[31:0] __l10_next[63:0];
	(*non_volatile*) reg[31:0] __l39_next[127:0];
	(*non_volatile*) reg[31:0] __l54_next;
	(*non_volatile*) reg[31:0] __l64_next[31:0];
	(*non_volatile*) reg signed[31:0] __l75_next;
	(*non_volatile*) reg[31:0] __l76_next;
	(*non_volatile*) reg signed[31:0] __l9_next;
	wire[31:0] __l10[63:0];
	assign __l10[0] = {__var[11]};
	assign __l10[1] = {__var[12]};
	assign __l10[2] = {__var[13]};
	assign __l10[3] = {__var[14]};
	assign __l10[4] = {__var[15]};
	assign __l10[5] = {__var[16]};
	assign __l10[6] = {__var[17]};
	assign __l10[7] = {__var[18]};
	assign __l10[8] = {__var[19]};
	assign __l10[9] = {__var[20]};
	assign __l10[10] = {__var[21]};
	assign __l10[11] = {__var[22]};
	assign __l10[12] = {__var[23]};
	assign __l10[13] = {__var[24]};
	assign __l10[14] = {__var[25]};
	assign __l10[15] = {__var[26]};
	assign __l10[16] = {__var[27]};
	assign __l10[17] = {__var[28]};
	assign __l10[18] = {__var[29]};
	assign __l10[19] = {__var[30]};
	assign __l10[20] = {__var[31]};
	assign __l10[21] = {__var[32]};
	assign __l10[22] = {__var[33]};
	assign __l10[23] = {__var[34]};
	assign __l10[24] = {__var[35]};
	assign __l10[25] = {__var[36]};
	assign __l10[26] = {__var[37]};
	assign __l10[27] = {__var[38]};
	assign __l10[28] = {__var[39]};
	assign __l10[29] = {__var[40]};
	assign __l10[30] = {__var[41]};
	assign __l10[31] = {__var[42]};
	assign __l10[32] = {__var[43]};
	assign __l10[33] = {__var[44]};
	assign __l10[34] = {__var[45]};
	assign __l10[35] = {__var[46]};
	assign __l10[36] = {__var[47]};
	assign __l10[37] = {__var[48]};
	assign __l10[38] = {__var[49]};
	assign __l10[39] = {__var[50]};
	assign __l10[40] = {__var[51]};
	assign __l10[41] = {__var[52]};
	assign __l10[42] = {__var[53]};
	assign __l10[43] = {__var[54]};
	assign __l10[44] = {__var[55]};
	assign __l10[45] = {__var[56]};
	assign __l10[46] = {__var[57]};
	assign __l10[47] = {__var[58]};
	assign __l10[48] = {__var[59]};
	assign __l10[49] = {__var[60]};
	assign __l10[50] = {__var[61]};
	assign __l10[51] = {__var[62]};
	assign __l10[52] = {__var[63]};
	assign __l10[53] = {__var[64]};
	assign __l10[54] = {__var[65]};
	assign __l10[55] = {__var[66]};
	assign __l10[56] = {__var[67]};
	assign __l10[57] = {__var[68]};
	assign __l10[58] = {__var[69]};
	assign __l10[59] = {__var[70]};
	assign __l10[60] = {__var[71]};
	assign __l10[61] = {__var[72]};
	assign __l10[62] = {__var[73]};
	assign __l10[63] = {__var[74]};
	wire[31:0] __l39[127:0];
	assign __l39[0] = {__var[75]};
	assign __l39[1] = {__var[76]};
	assign __l39[2] = {__var[77]};
	assign __l39[3] = {__var[78]};
	assign __l39[4] = {__var[79]};
	assign __l39[5] = {__var[80]};
	assign __l39[6] = {__var[81]};
	assign __l39[7] = {__var[82]};
	assign __l39[8] = {__var[83]};
	assign __l39[9] = {__var[84]};
	assign __l39[10] = {__var[85]};
	assign __l39[11] = {__var[86]};
	assign __l39[12] = {__var[87]};
	assign __l39[13] = {__var[88]};
	assign __l39[14] = {__var[89]};
	assign __l39[15] = {__var[90]};
	assign __l39[16] = {__var[91]};
	assign __l39[17] = {__var[92]};
	assign __l39[18] = {__var[93]};
	assign __l39[19] = {__var[94]};
	assign __l39[20] = {__var[95]};
	assign __l39[21] = {__var[96]};
	assign __l39[22] = {__var[97]};
	assign __l39[23] = {__var[98]};
	assign __l39[24] = {__var[99]};
	assign __l39[25] = {__var[100]};
	assign __l39[26] = {__var[101]};
	assign __l39[27] = {__var[102]};
	assign __l39[28] = {__var[103]};
	assign __l39[29] = {__var[104]};
	assign __l39[30] = {__var[105]};
	assign __l39[31] = {__var[106]};
	assign __l39[32] = {__var[107]};
	assign __l39[33] = {__var[108]};
	assign __l39[34] = {__var[109]};
	assign __l39[35] = {__var[110]};
	assign __l39[36] = {__var[111]};
	assign __l39[37] = {__var[112]};
	assign __l39[38] = {__var[113]};
	assign __l39[39] = {__var[114]};
	assign __l39[40] = {__var[115]};
	assign __l39[41] = {__var[116]};
	assign __l39[42] = {__var[117]};
	assign __l39[43] = {__var[118]};
	assign __l39[44] = {__var[119]};
	assign __l39[45] = {__var[120]};
	assign __l39[46] = {__var[121]};
	assign __l39[47] = {__var[122]};
	assign __l39[48] = {__var[123]};
	assign __l39[49] = {__var[124]};
	assign __l39[50] = {__var[125]};
	assign __l39[51] = {__var[126]};
	assign __l39[52] = {__var[127]};
	assign __l39[53] = {__var[128]};
	assign __l39[54] = {__var[129]};
	assign __l39[55] = {__var[130]};
	assign __l39[56] = {__var[131]};
	assign __l39[57] = {__var[132]};
	assign __l39[58] = {__var[133]};
	assign __l39[59] = {__var[134]};
	assign __l39[60] = {__var[135]};
	assign __l39[61] = {__var[136]};
	assign __l39[62] = {__var[137]};
	assign __l39[63] = {__var[138]};
	assign __l39[64] = {__var[139]};
	assign __l39[65] = {__var[140]};
	assign __l39[66] = {__var[141]};
	assign __l39[67] = {__var[142]};
	assign __l39[68] = {__var[143]};
	assign __l39[69] = {__var[144]};
	assign __l39[70] = {__var[145]};
	assign __l39[71] = {__var[146]};
	assign __l39[72] = {__var[147]};
	assign __l39[73] = {__var[148]};
	assign __l39[74] = {__var[149]};
	assign __l39[75] = {__var[150]};
	assign __l39[76] = {__var[151]};
	assign __l39[77] = {__var[152]};
	assign __l39[78] = {__var[153]};
	assign __l39[79] = {__var[154]};
	assign __l39[80] = {__var[155]};
	assign __l39[81] = {__var[156]};
	assign __l39[82] = {__var[157]};
	assign __l39[83] = {__var[158]};
	assign __l39[84] = {__var[159]};
	assign __l39[85] = {__var[160]};
	assign __l39[86] = {__var[161]};
	assign __l39[87] = {__var[162]};
	assign __l39[88] = {__var[163]};
	assign __l39[89] = {__var[164]};
	assign __l39[90] = {__var[165]};
	assign __l39[91] = {__var[166]};
	assign __l39[92] = {__var[167]};
	assign __l39[93] = {__var[168]};
	assign __l39[94] = {__var[169]};
	assign __l39[95] = {__var[170]};
	assign __l39[96] = {__var[171]};
	assign __l39[97] = {__var[172]};
	assign __l39[98] = {__var[173]};
	assign __l39[99] = {__var[174]};
	assign __l39[100] = {__var[175]};
	assign __l39[101] = {__var[176]};
	assign __l39[102] = {__var[177]};
	assign __l39[103] = {__var[178]};
	assign __l39[104] = {__var[179]};
	assign __l39[105] = {__var[180]};
	assign __l39[106] = {__var[181]};
	assign __l39[107] = {__var[182]};
	assign __l39[108] = {__var[183]};
	assign __l39[109] = {__var[184]};
	assign __l39[110] = {__var[185]};
	assign __l39[111] = {__var[186]};
	assign __l39[112] = {__var[187]};
	assign __l39[113] = {__var[188]};
	assign __l39[114] = {__var[189]};
	assign __l39[115] = {__var[190]};
	assign __l39[116] = {__var[191]};
	assign __l39[117] = {__var[192]};
	assign __l39[118] = {__var[193]};
	assign __l39[119] = {__var[194]};
	assign __l39[120] = {__var[195]};
	assign __l39[121] = {__var[196]};
	assign __l39[122] = {__var[197]};
	assign __l39[123] = {__var[198]};
	assign __l39[124] = {__var[199]};
	assign __l39[125] = {__var[200]};
	assign __l39[126] = {__var[201]};
	assign __l39[127] = {__var[202]};
	wire[31:0] __l54;
	assign __l54 = {__var[203]};
	wire[31:0] __l64[31:0];
	assign __l64[0] = {__var[204]};
	assign __l64[1] = {__var[205]};
	assign __l64[2] = {__var[206]};
	assign __l64[3] = {__var[207]};
	assign __l64[4] = {__var[208]};
	assign __l64[5] = {__var[209]};
	assign __l64[6] = {__var[210]};
	assign __l64[7] = {__var[211]};
	assign __l64[8] = {__var[212]};
	assign __l64[9] = {__var[213]};
	assign __l64[10] = {__var[214]};
	assign __l64[11] = {__var[215]};
	assign __l64[12] = {__var[216]};
	assign __l64[13] = {__var[217]};
	assign __l64[14] = {__var[218]};
	assign __l64[15] = {__var[219]};
	assign __l64[16] = {__var[220]};
	assign __l64[17] = {__var[221]};
	assign __l64[18] = {__var[222]};
	assign __l64[19] = {__var[223]};
	assign __l64[20] = {__var[224]};
	assign __l64[21] = {__var[225]};
	assign __l64[22] = {__var[226]};
	assign __l64[23] = {__var[227]};
	assign __l64[24] = {__var[228]};
	assign __l64[25] = {__var[229]};
	assign __l64[26] = {__var[230]};
	assign __l64[27] = {__var[231]};
	assign __l64[28] = {__var[232]};
	assign __l64[29] = {__var[233]};
	assign __l64[30] = {__var[234]};
	assign __l64[31] = {__var[235]};
	wire signed[31:0] __l75;
	assign __l75 = {__var[236]};
	wire[31:0] __l76;
	assign __l76 = {__var[237]};
	wire signed[31:0] __l9;
	assign __l9 = {__var[10]};
	wire __x1;
	assign __x1 = {__var[9]};
	reg[238:0] __update_queue;
	wire __there_are_updates;
	wire __apply_updates;
	wire __there_were_tasks;
	wire __all_final;
	wire __continue;
	wire __reset;
	reg __x1_prev;
	wire __x1_posedge;
	wire __any_triggers;
	reg[31:0] __open_loop = 0;
	wire __open_loop_tick;
	wire[31:0] __l11;
	wire[31:0] __l13;
	wire[31:0] __l14;
	(*non_volatile*) reg[31:0] __l15;
	wire __l16;
	(*non_volatile*) reg[3:0] __l18;
	wire[31:0] __l24;
	(*non_volatile*) reg __l26;
	(*non_volatile*) reg[1:0] __l27;
	(*non_volatile*) reg __l28;
	(*non_volatile*) reg __l30;
	(*non_volatile*) reg __l31;
	(*non_volatile*) reg __l32;
	(*non_volatile*) reg __l33;
	(*non_volatile*) reg __l34;
	wire[6:0] __l40;
	wire[6:0] __l41;
	wire[31:0] __l42;
	wire[31:0] __l43;
	wire[6:0] __l44;
	wire[31:0] __l47;
	wire[31:0] __l50;
	wire[31:0] __l55;
	wire[31:0] __l56;
	wire[31:0] __l60;
	wire[31:0] __l67;
	wire[31:0] __l68;
	wire[4:0] __l69;
	assign __l11 = __l10[__l56];
	assign __l55 = (__l54 + 4);
	assign __l56 = (__l54 >> 2);
	assign __l47 = {(__l11[15] ? 16'b0000000000000001 : 16'b0000000000000000),__l11[15:0]};
	assign __l50 = {__l55[31:28],__l11[25:0],2'b00};
	assign __l24 = (__l55 + (__l47 << 2));
	assign __l67 = __l64[__l11[25:21]];
	assign __l68 = __l64[__l11[20:16]];
	assign __l69 = (__l33 ? __l11[15:11] : __l11[20:16]);
	assign __l16 = (__l15 == 32'b00000000000000000000000000000000);
	assign __l13 = (__l27[1] ? __l68 : __l67);
	assign __l14 = (__l27[1] ? (__l27[0] ? __l67 : __l11[10:6]) : (__l27[0] ? __l47 : __l68));
	assign __l42 = __l39[__l40];
	assign __l43 = __l39[__l41];
	assign __l40 = (__l15 >> 2);
	assign __l44 = (__l15 >> 2);
	assign __l60 = (__l31 ? __l42 : __l15);
	always @(__l13 or __l14 or __l18) begin
		case (__l18)
			4'b0000: __l15 = (__l13 << __l14);
			4'b0001: __l15 = (__l13 >> __l14);
			4'b0010: __l15 = (__l13 >>> __l14);
			4'b0011: __l15 = (__l13 + __l14);
			4'b0100: __l15 = (__l13 - __l14);
			4'b0101: __l15 = (__l13 & __l14);
			4'b0110: __l15 = (__l13 | __l14);
			4'b0111: __l15 = (__l13 ^ __l14);
			4'b1000: __l15 = (!(__l13 | __l14));
			4'b1001: __l15 = ((__l13 < __l14) ? 1 : 0);
			4'b1010: __l15 = (__l14 << 16);
			default: __l15 = 0;
		endcase
	end 
	always @(__l11 or __l26) begin
		if ((__l26 == 0)) begin
			case (__l11[31:26])
				6'd4: __l18 = 4'b0100;
				6'd8: __l18 = 4'b0011;
				6'd10: __l18 = 4'b1001;
				6'd12: __l18 = 4'b0101;
				6'd13: __l18 = 4'b0110;
				6'd14: __l18 = 4'b0111;
				6'd15: __l18 = 4'b1010;
				6'd35: __l18 = 4'b0011;
				6'd43: __l18 = 4'b0011;
				default: __l18 = 0;
			endcase
		end 
		else begin
			case (__l11[5:0])
				6'd0: __l18 = 4'b0000;
				6'd2: __l18 = 4'b0001;
				6'd3: __l18 = 4'b0010;
				6'd6: __l18 = 4'b0001;
				6'd7: __l18 = 4'b0010;
				6'd32: __l18 = 4'b0011;
				6'd34: __l18 = 4'b0100;
				6'd36: __l18 = 4'b0101;
				6'd37: __l18 = 4'b0110;
				6'd38: __l18 = 4'b0111;
				6'd39: __l18 = 4'b1000;
				6'd42: __l18 = 4'b1001;
				default: __l18 = 0;
			endcase
		end 
	end 
	always @(__l11) begin
		case (__l11[31:26])
			6'd0: if ((__l11[5:0] == 6'd13)) begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b00;
				__l34 = 0;
			end 
			else 
				if ((__l11[5:0] < 6'd4)) begin
					__l33 = 1;
					__l30 = 0;
					__l28 = 0;
					__l31 = 0;
					__l26 = 1;
					__l32 = 0;
					__l27 = 2'b10;
					__l34 = 1;
				end 
				else 
					if ((__l11[5:0] < 6'd8)) begin
						__l33 = 1;
						__l30 = 0;
						__l28 = 0;
						__l31 = 0;
						__l26 = 1;
						__l32 = 0;
						__l27 = 2'b11;
						__l34 = 1;
					end 
					else begin
						__l33 = 1;
						__l30 = 0;
						__l28 = 0;
						__l31 = 0;
						__l26 = 1;
						__l32 = 0;
						__l27 = 2'b00;
						__l34 = 1;
					end 
			6'd2: begin
				__l33 = 0;
				__l30 = 1;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b00;
				__l34 = 0;
			end 
			6'd4: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 1;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b00;
				__l34 = 0;
			end 
			6'd8: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd10: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd12: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd13: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd14: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd15: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd35: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 1;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b01;
				__l34 = 1;
			end 
			6'd43: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 1;
				__l27 = 2'b01;
				__l34 = 0;
			end 
			default: begin
				__l33 = 0;
				__l30 = 0;
				__l28 = 0;
				__l31 = 0;
				__l26 = 0;
				__l32 = 0;
				__l27 = 2'b00;
				__l34 = 0;
			end 
		endcase
	end 
	reg[15:0] __task_id[0:0];
	reg[15:0] __state[0:0];
	reg[15:0] __paused[0:0];
	always @(posedge __clk) begin : __buf_block
		__read_buf[3] <= ((__in_valid && __in_read) << __in_vid);
		__read_buf[2] <= __read_buf[3];
		__write_buf[3] <= ((__in_valid && (!__in_read)) << __in_vid);
		__write_buf[2] <= __write_buf[3];
		__in_buf[3] <= __in_data;
		__in_buf[2] <= __in_buf[3];
	end 
	assign __read = __read_buf[2];
	assign __write = __write_buf[2];
	assign __in = __in_buf[2];
	assign __there_are_updates = (|__update_queue);
	assign __apply_updates = (__read[1] || __open_loop_tick);
	assign __there_were_tasks = (|{(__task_id[0] != 0)});
	assign __all_final = (&{(__state[0] == 5)});
	assign __continue = __read[3];
	assign __reset = __read[4];
	always @(posedge __clk) begin
		__x1_prev <= __x1;
	end 
	assign __x1_posedge = ((__x1_prev == 0) && (__x1 == 1));
	assign __any_triggers = (|{__x1_posedge});
	always @(posedge __clk) __open_loop <= (__read[5] ? __in : (__open_loop_tick ? (__open_loop - 1) : __open_loop));
	assign __open_loop_tick = (__all_final && ((!__any_triggers) && (__open_loop > 0)));
	always @(posedge __clk) begin
		__state[0] = (__x1_posedge ? 0 : __state[0]);
		if (((__state[0] == 0) && (!__paused[0]))) begin
			if (__l34) begin
				__l64_next[__l69] <= __l60;
				__update_queue[(204 + (__l69 * 1))+:1] <= (~0);
			end 
			if (__l32) begin
				__l39_next[__l44] <= __l68;
				__update_queue[(75 + (__l44 * 1))+:1] <= (~0);
			end 
			if ((__l11[5:0] == 6'd13)) 
				__state[0] = 1;
			else 
				__state[0] = 4;
		end 
		if (((__state[0] == 1) && (!__paused[0]))) begin
			__paused[0] = 1;
			__task_id[0] = 1;
			__state[0] = 2;
		end 
		if (((__state[0] == 2) && (!__paused[0]))) begin
			__paused[0] = 1;
			__task_id[0] = 2;
			__state[0] = 3;
		end 
		if (((__state[0] == 3) && (!__paused[0]))) begin
			__paused[0] = 1;
			__task_id[0] = 3;
			__state[0] = 4;
		end 
		if (((__state[0] == 4) && (!__paused[0]))) begin
			if (__l30) begin
				__l54_next <= __l50;
				__update_queue[203+:1] <= (~0);
			end 
			else 
				if ((__l28 & __l16)) begin
					__l54_next <= __l24;
					__update_queue[203+:1] <= (~0);
				end 
				else begin
					__l54_next <= __l55;
					__update_queue[203+:1] <= (~0);
				end 
			__state[0] = 5;
		end 
		if (((__state[0] == 5) && (!__paused[0]))) begin
			__state[0] = 5;
		end 
		__paused[0] = (__reset ? 1 : (__continue ? 0 : __paused[0]));
		__task_id[0] = (__reset ? 65535 : (__continue ? 0 : __task_id[0]));
		__state[0] = (__reset ? 5 : __state[0]);
		__var[9][0:0] <= (__open_loop_tick ? (~__x1) : (__read[9] ? __in : __var[9]));
		__var[10][31:0] <= (__read[10] ? __in : ((__apply_updates && __update_queue[10]) ? __l9_next[31:0] : __var[10]));
		__var[11][31:0] <= (__read[11] ? __in : ((__apply_updates && __update_queue[11]) ? __l10_next[0][31:0] : __var[11]));
		__var[12][31:0] <= (__read[12] ? __in : ((__apply_updates && __update_queue[12]) ? __l10_next[1][31:0] : __var[12]));
		__var[13][31:0] <= (__read[13] ? __in : ((__apply_updates && __update_queue[13]) ? __l10_next[2][31:0] : __var[13]));
		__var[14][31:0] <= (__read[14] ? __in : ((__apply_updates && __update_queue[14]) ? __l10_next[3][31:0] : __var[14]));
		__var[15][31:0] <= (__read[15] ? __in : ((__apply_updates && __update_queue[15]) ? __l10_next[4][31:0] : __var[15]));
		__var[16][31:0] <= (__read[16] ? __in : ((__apply_updates && __update_queue[16]) ? __l10_next[5][31:0] : __var[16]));
		__var[17][31:0] <= (__read[17] ? __in : ((__apply_updates && __update_queue[17]) ? __l10_next[6][31:0] : __var[17]));
		__var[18][31:0] <= (__read[18] ? __in : ((__apply_updates && __update_queue[18]) ? __l10_next[7][31:0] : __var[18]));
		__var[19][31:0] <= (__read[19] ? __in : ((__apply_updates && __update_queue[19]) ? __l10_next[8][31:0] : __var[19]));
		__var[20][31:0] <= (__read[20] ? __in : ((__apply_updates && __update_queue[20]) ? __l10_next[9][31:0] : __var[20]));
		__var[21][31:0] <= (__read[21] ? __in : ((__apply_updates && __update_queue[21]) ? __l10_next[10][31:0] : __var[21]));
		__var[22][31:0] <= (__read[22] ? __in : ((__apply_updates && __update_queue[22]) ? __l10_next[11][31:0] : __var[22]));
		__var[23][31:0] <= (__read[23] ? __in : ((__apply_updates && __update_queue[23]) ? __l10_next[12][31:0] : __var[23]));
		__var[24][31:0] <= (__read[24] ? __in : ((__apply_updates && __update_queue[24]) ? __l10_next[13][31:0] : __var[24]));
		__var[25][31:0] <= (__read[25] ? __in : ((__apply_updates && __update_queue[25]) ? __l10_next[14][31:0] : __var[25]));
		__var[26][31:0] <= (__read[26] ? __in : ((__apply_updates && __update_queue[26]) ? __l10_next[15][31:0] : __var[26]));
		__var[27][31:0] <= (__read[27] ? __in : ((__apply_updates && __update_queue[27]) ? __l10_next[16][31:0] : __var[27]));
		__var[28][31:0] <= (__read[28] ? __in : ((__apply_updates && __update_queue[28]) ? __l10_next[17][31:0] : __var[28]));
		__var[29][31:0] <= (__read[29] ? __in : ((__apply_updates && __update_queue[29]) ? __l10_next[18][31:0] : __var[29]));
		__var[30][31:0] <= (__read[30] ? __in : ((__apply_updates && __update_queue[30]) ? __l10_next[19][31:0] : __var[30]));
		__var[31][31:0] <= (__read[31] ? __in : ((__apply_updates && __update_queue[31]) ? __l10_next[20][31:0] : __var[31]));
		__var[32][31:0] <= (__read[32] ? __in : ((__apply_updates && __update_queue[32]) ? __l10_next[21][31:0] : __var[32]));
		__var[33][31:0] <= (__read[33] ? __in : ((__apply_updates && __update_queue[33]) ? __l10_next[22][31:0] : __var[33]));
		__var[34][31:0] <= (__read[34] ? __in : ((__apply_updates && __update_queue[34]) ? __l10_next[23][31:0] : __var[34]));
		__var[35][31:0] <= (__read[35] ? __in : ((__apply_updates && __update_queue[35]) ? __l10_next[24][31:0] : __var[35]));
		__var[36][31:0] <= (__read[36] ? __in : ((__apply_updates && __update_queue[36]) ? __l10_next[25][31:0] : __var[36]));
		__var[37][31:0] <= (__read[37] ? __in : ((__apply_updates && __update_queue[37]) ? __l10_next[26][31:0] : __var[37]));
		__var[38][31:0] <= (__read[38] ? __in : ((__apply_updates && __update_queue[38]) ? __l10_next[27][31:0] : __var[38]));
		__var[39][31:0] <= (__read[39] ? __in : ((__apply_updates && __update_queue[39]) ? __l10_next[28][31:0] : __var[39]));
		__var[40][31:0] <= (__read[40] ? __in : ((__apply_updates && __update_queue[40]) ? __l10_next[29][31:0] : __var[40]));
		__var[41][31:0] <= (__read[41] ? __in : ((__apply_updates && __update_queue[41]) ? __l10_next[30][31:0] : __var[41]));
		__var[42][31:0] <= (__read[42] ? __in : ((__apply_updates && __update_queue[42]) ? __l10_next[31][31:0] : __var[42]));
		__var[43][31:0] <= (__read[43] ? __in : ((__apply_updates && __update_queue[43]) ? __l10_next[32][31:0] : __var[43]));
		__var[44][31:0] <= (__read[44] ? __in : ((__apply_updates && __update_queue[44]) ? __l10_next[33][31:0] : __var[44]));
		__var[45][31:0] <= (__read[45] ? __in : ((__apply_updates && __update_queue[45]) ? __l10_next[34][31:0] : __var[45]));
		__var[46][31:0] <= (__read[46] ? __in : ((__apply_updates && __update_queue[46]) ? __l10_next[35][31:0] : __var[46]));
		__var[47][31:0] <= (__read[47] ? __in : ((__apply_updates && __update_queue[47]) ? __l10_next[36][31:0] : __var[47]));
		__var[48][31:0] <= (__read[48] ? __in : ((__apply_updates && __update_queue[48]) ? __l10_next[37][31:0] : __var[48]));
		__var[49][31:0] <= (__read[49] ? __in : ((__apply_updates && __update_queue[49]) ? __l10_next[38][31:0] : __var[49]));
		__var[50][31:0] <= (__read[50] ? __in : ((__apply_updates && __update_queue[50]) ? __l10_next[39][31:0] : __var[50]));
		__var[51][31:0] <= (__read[51] ? __in : ((__apply_updates && __update_queue[51]) ? __l10_next[40][31:0] : __var[51]));
		__var[52][31:0] <= (__read[52] ? __in : ((__apply_updates && __update_queue[52]) ? __l10_next[41][31:0] : __var[52]));
		__var[53][31:0] <= (__read[53] ? __in : ((__apply_updates && __update_queue[53]) ? __l10_next[42][31:0] : __var[53]));
		__var[54][31:0] <= (__read[54] ? __in : ((__apply_updates && __update_queue[54]) ? __l10_next[43][31:0] : __var[54]));
		__var[55][31:0] <= (__read[55] ? __in : ((__apply_updates && __update_queue[55]) ? __l10_next[44][31:0] : __var[55]));
		__var[56][31:0] <= (__read[56] ? __in : ((__apply_updates && __update_queue[56]) ? __l10_next[45][31:0] : __var[56]));
		__var[57][31:0] <= (__read[57] ? __in : ((__apply_updates && __update_queue[57]) ? __l10_next[46][31:0] : __var[57]));
		__var[58][31:0] <= (__read[58] ? __in : ((__apply_updates && __update_queue[58]) ? __l10_next[47][31:0] : __var[58]));
		__var[59][31:0] <= (__read[59] ? __in : ((__apply_updates && __update_queue[59]) ? __l10_next[48][31:0] : __var[59]));
		__var[60][31:0] <= (__read[60] ? __in : ((__apply_updates && __update_queue[60]) ? __l10_next[49][31:0] : __var[60]));
		__var[61][31:0] <= (__read[61] ? __in : ((__apply_updates && __update_queue[61]) ? __l10_next[50][31:0] : __var[61]));
		__var[62][31:0] <= (__read[62] ? __in : ((__apply_updates && __update_queue[62]) ? __l10_next[51][31:0] : __var[62]));
		__var[63][31:0] <= (__read[63] ? __in : ((__apply_updates && __update_queue[63]) ? __l10_next[52][31:0] : __var[63]));
		__var[64][31:0] <= (__read[64] ? __in : ((__apply_updates && __update_queue[64]) ? __l10_next[53][31:0] : __var[64]));
		__var[65][31:0] <= (__read[65] ? __in : ((__apply_updates && __update_queue[65]) ? __l10_next[54][31:0] : __var[65]));
		__var[66][31:0] <= (__read[66] ? __in : ((__apply_updates && __update_queue[66]) ? __l10_next[55][31:0] : __var[66]));
		__var[67][31:0] <= (__read[67] ? __in : ((__apply_updates && __update_queue[67]) ? __l10_next[56][31:0] : __var[67]));
		__var[68][31:0] <= (__read[68] ? __in : ((__apply_updates && __update_queue[68]) ? __l10_next[57][31:0] : __var[68]));
		__var[69][31:0] <= (__read[69] ? __in : ((__apply_updates && __update_queue[69]) ? __l10_next[58][31:0] : __var[69]));
		__var[70][31:0] <= (__read[70] ? __in : ((__apply_updates && __update_queue[70]) ? __l10_next[59][31:0] : __var[70]));
		__var[71][31:0] <= (__read[71] ? __in : ((__apply_updates && __update_queue[71]) ? __l10_next[60][31:0] : __var[71]));
		__var[72][31:0] <= (__read[72] ? __in : ((__apply_updates && __update_queue[72]) ? __l10_next[61][31:0] : __var[72]));
		__var[73][31:0] <= (__read[73] ? __in : ((__apply_updates && __update_queue[73]) ? __l10_next[62][31:0] : __var[73]));
		__var[74][31:0] <= (__read[74] ? __in : ((__apply_updates && __update_queue[74]) ? __l10_next[63][31:0] : __var[74]));
		__var[75][31:0] <= (__read[75] ? __in : ((__apply_updates && __update_queue[75]) ? __l39_next[0][31:0] : __var[75]));
		__var[76][31:0] <= (__read[76] ? __in : ((__apply_updates && __update_queue[76]) ? __l39_next[1][31:0] : __var[76]));
		__var[77][31:0] <= (__read[77] ? __in : ((__apply_updates && __update_queue[77]) ? __l39_next[2][31:0] : __var[77]));
		__var[78][31:0] <= (__read[78] ? __in : ((__apply_updates && __update_queue[78]) ? __l39_next[3][31:0] : __var[78]));
		__var[79][31:0] <= (__read[79] ? __in : ((__apply_updates && __update_queue[79]) ? __l39_next[4][31:0] : __var[79]));
		__var[80][31:0] <= (__read[80] ? __in : ((__apply_updates && __update_queue[80]) ? __l39_next[5][31:0] : __var[80]));
		__var[81][31:0] <= (__read[81] ? __in : ((__apply_updates && __update_queue[81]) ? __l39_next[6][31:0] : __var[81]));
		__var[82][31:0] <= (__read[82] ? __in : ((__apply_updates && __update_queue[82]) ? __l39_next[7][31:0] : __var[82]));
		__var[83][31:0] <= (__read[83] ? __in : ((__apply_updates && __update_queue[83]) ? __l39_next[8][31:0] : __var[83]));
		__var[84][31:0] <= (__read[84] ? __in : ((__apply_updates && __update_queue[84]) ? __l39_next[9][31:0] : __var[84]));
		__var[85][31:0] <= (__read[85] ? __in : ((__apply_updates && __update_queue[85]) ? __l39_next[10][31:0] : __var[85]));
		__var[86][31:0] <= (__read[86] ? __in : ((__apply_updates && __update_queue[86]) ? __l39_next[11][31:0] : __var[86]));
		__var[87][31:0] <= (__read[87] ? __in : ((__apply_updates && __update_queue[87]) ? __l39_next[12][31:0] : __var[87]));
		__var[88][31:0] <= (__read[88] ? __in : ((__apply_updates && __update_queue[88]) ? __l39_next[13][31:0] : __var[88]));
		__var[89][31:0] <= (__read[89] ? __in : ((__apply_updates && __update_queue[89]) ? __l39_next[14][31:0] : __var[89]));
		__var[90][31:0] <= (__read[90] ? __in : ((__apply_updates && __update_queue[90]) ? __l39_next[15][31:0] : __var[90]));
		__var[91][31:0] <= (__read[91] ? __in : ((__apply_updates && __update_queue[91]) ? __l39_next[16][31:0] : __var[91]));
		__var[92][31:0] <= (__read[92] ? __in : ((__apply_updates && __update_queue[92]) ? __l39_next[17][31:0] : __var[92]));
		__var[93][31:0] <= (__read[93] ? __in : ((__apply_updates && __update_queue[93]) ? __l39_next[18][31:0] : __var[93]));
		__var[94][31:0] <= (__read[94] ? __in : ((__apply_updates && __update_queue[94]) ? __l39_next[19][31:0] : __var[94]));
		__var[95][31:0] <= (__read[95] ? __in : ((__apply_updates && __update_queue[95]) ? __l39_next[20][31:0] : __var[95]));
		__var[96][31:0] <= (__read[96] ? __in : ((__apply_updates && __update_queue[96]) ? __l39_next[21][31:0] : __var[96]));
		__var[97][31:0] <= (__read[97] ? __in : ((__apply_updates && __update_queue[97]) ? __l39_next[22][31:0] : __var[97]));
		__var[98][31:0] <= (__read[98] ? __in : ((__apply_updates && __update_queue[98]) ? __l39_next[23][31:0] : __var[98]));
		__var[99][31:0] <= (__read[99] ? __in : ((__apply_updates && __update_queue[99]) ? __l39_next[24][31:0] : __var[99]));
		__var[100][31:0] <= (__read[100] ? __in : ((__apply_updates && __update_queue[100]) ? __l39_next[25][31:0] : __var[100]));
		__var[101][31:0] <= (__read[101] ? __in : ((__apply_updates && __update_queue[101]) ? __l39_next[26][31:0] : __var[101]));
		__var[102][31:0] <= (__read[102] ? __in : ((__apply_updates && __update_queue[102]) ? __l39_next[27][31:0] : __var[102]));
		__var[103][31:0] <= (__read[103] ? __in : ((__apply_updates && __update_queue[103]) ? __l39_next[28][31:0] : __var[103]));
		__var[104][31:0] <= (__read[104] ? __in : ((__apply_updates && __update_queue[104]) ? __l39_next[29][31:0] : __var[104]));
		__var[105][31:0] <= (__read[105] ? __in : ((__apply_updates && __update_queue[105]) ? __l39_next[30][31:0] : __var[105]));
		__var[106][31:0] <= (__read[106] ? __in : ((__apply_updates && __update_queue[106]) ? __l39_next[31][31:0] : __var[106]));
		__var[107][31:0] <= (__read[107] ? __in : ((__apply_updates && __update_queue[107]) ? __l39_next[32][31:0] : __var[107]));
		__var[108][31:0] <= (__read[108] ? __in : ((__apply_updates && __update_queue[108]) ? __l39_next[33][31:0] : __var[108]));
		__var[109][31:0] <= (__read[109] ? __in : ((__apply_updates && __update_queue[109]) ? __l39_next[34][31:0] : __var[109]));
		__var[110][31:0] <= (__read[110] ? __in : ((__apply_updates && __update_queue[110]) ? __l39_next[35][31:0] : __var[110]));
		__var[111][31:0] <= (__read[111] ? __in : ((__apply_updates && __update_queue[111]) ? __l39_next[36][31:0] : __var[111]));
		__var[112][31:0] <= (__read[112] ? __in : ((__apply_updates && __update_queue[112]) ? __l39_next[37][31:0] : __var[112]));
		__var[113][31:0] <= (__read[113] ? __in : ((__apply_updates && __update_queue[113]) ? __l39_next[38][31:0] : __var[113]));
		__var[114][31:0] <= (__read[114] ? __in : ((__apply_updates && __update_queue[114]) ? __l39_next[39][31:0] : __var[114]));
		__var[115][31:0] <= (__read[115] ? __in : ((__apply_updates && __update_queue[115]) ? __l39_next[40][31:0] : __var[115]));
		__var[116][31:0] <= (__read[116] ? __in : ((__apply_updates && __update_queue[116]) ? __l39_next[41][31:0] : __var[116]));
		__var[117][31:0] <= (__read[117] ? __in : ((__apply_updates && __update_queue[117]) ? __l39_next[42][31:0] : __var[117]));
		__var[118][31:0] <= (__read[118] ? __in : ((__apply_updates && __update_queue[118]) ? __l39_next[43][31:0] : __var[118]));
		__var[119][31:0] <= (__read[119] ? __in : ((__apply_updates && __update_queue[119]) ? __l39_next[44][31:0] : __var[119]));
		__var[120][31:0] <= (__read[120] ? __in : ((__apply_updates && __update_queue[120]) ? __l39_next[45][31:0] : __var[120]));
		__var[121][31:0] <= (__read[121] ? __in : ((__apply_updates && __update_queue[121]) ? __l39_next[46][31:0] : __var[121]));
		__var[122][31:0] <= (__read[122] ? __in : ((__apply_updates && __update_queue[122]) ? __l39_next[47][31:0] : __var[122]));
		__var[123][31:0] <= (__read[123] ? __in : ((__apply_updates && __update_queue[123]) ? __l39_next[48][31:0] : __var[123]));
		__var[124][31:0] <= (__read[124] ? __in : ((__apply_updates && __update_queue[124]) ? __l39_next[49][31:0] : __var[124]));
		__var[125][31:0] <= (__read[125] ? __in : ((__apply_updates && __update_queue[125]) ? __l39_next[50][31:0] : __var[125]));
		__var[126][31:0] <= (__read[126] ? __in : ((__apply_updates && __update_queue[126]) ? __l39_next[51][31:0] : __var[126]));
		__var[127][31:0] <= (__read[127] ? __in : ((__apply_updates && __update_queue[127]) ? __l39_next[52][31:0] : __var[127]));
		__var[128][31:0] <= (__read[128] ? __in : ((__apply_updates && __update_queue[128]) ? __l39_next[53][31:0] : __var[128]));
		__var[129][31:0] <= (__read[129] ? __in : ((__apply_updates && __update_queue[129]) ? __l39_next[54][31:0] : __var[129]));
		__var[130][31:0] <= (__read[130] ? __in : ((__apply_updates && __update_queue[130]) ? __l39_next[55][31:0] : __var[130]));
		__var[131][31:0] <= (__read[131] ? __in : ((__apply_updates && __update_queue[131]) ? __l39_next[56][31:0] : __var[131]));
		__var[132][31:0] <= (__read[132] ? __in : ((__apply_updates && __update_queue[132]) ? __l39_next[57][31:0] : __var[132]));
		__var[133][31:0] <= (__read[133] ? __in : ((__apply_updates && __update_queue[133]) ? __l39_next[58][31:0] : __var[133]));
		__var[134][31:0] <= (__read[134] ? __in : ((__apply_updates && __update_queue[134]) ? __l39_next[59][31:0] : __var[134]));
		__var[135][31:0] <= (__read[135] ? __in : ((__apply_updates && __update_queue[135]) ? __l39_next[60][31:0] : __var[135]));
		__var[136][31:0] <= (__read[136] ? __in : ((__apply_updates && __update_queue[136]) ? __l39_next[61][31:0] : __var[136]));
		__var[137][31:0] <= (__read[137] ? __in : ((__apply_updates && __update_queue[137]) ? __l39_next[62][31:0] : __var[137]));
		__var[138][31:0] <= (__read[138] ? __in : ((__apply_updates && __update_queue[138]) ? __l39_next[63][31:0] : __var[138]));
		__var[139][31:0] <= (__read[139] ? __in : ((__apply_updates && __update_queue[139]) ? __l39_next[64][31:0] : __var[139]));
		__var[140][31:0] <= (__read[140] ? __in : ((__apply_updates && __update_queue[140]) ? __l39_next[65][31:0] : __var[140]));
		__var[141][31:0] <= (__read[141] ? __in : ((__apply_updates && __update_queue[141]) ? __l39_next[66][31:0] : __var[141]));
		__var[142][31:0] <= (__read[142] ? __in : ((__apply_updates && __update_queue[142]) ? __l39_next[67][31:0] : __var[142]));
		__var[143][31:0] <= (__read[143] ? __in : ((__apply_updates && __update_queue[143]) ? __l39_next[68][31:0] : __var[143]));
		__var[144][31:0] <= (__read[144] ? __in : ((__apply_updates && __update_queue[144]) ? __l39_next[69][31:0] : __var[144]));
		__var[145][31:0] <= (__read[145] ? __in : ((__apply_updates && __update_queue[145]) ? __l39_next[70][31:0] : __var[145]));
		__var[146][31:0] <= (__read[146] ? __in : ((__apply_updates && __update_queue[146]) ? __l39_next[71][31:0] : __var[146]));
		__var[147][31:0] <= (__read[147] ? __in : ((__apply_updates && __update_queue[147]) ? __l39_next[72][31:0] : __var[147]));
		__var[148][31:0] <= (__read[148] ? __in : ((__apply_updates && __update_queue[148]) ? __l39_next[73][31:0] : __var[148]));
		__var[149][31:0] <= (__read[149] ? __in : ((__apply_updates && __update_queue[149]) ? __l39_next[74][31:0] : __var[149]));
		__var[150][31:0] <= (__read[150] ? __in : ((__apply_updates && __update_queue[150]) ? __l39_next[75][31:0] : __var[150]));
		__var[151][31:0] <= (__read[151] ? __in : ((__apply_updates && __update_queue[151]) ? __l39_next[76][31:0] : __var[151]));
		__var[152][31:0] <= (__read[152] ? __in : ((__apply_updates && __update_queue[152]) ? __l39_next[77][31:0] : __var[152]));
		__var[153][31:0] <= (__read[153] ? __in : ((__apply_updates && __update_queue[153]) ? __l39_next[78][31:0] : __var[153]));
		__var[154][31:0] <= (__read[154] ? __in : ((__apply_updates && __update_queue[154]) ? __l39_next[79][31:0] : __var[154]));
		__var[155][31:0] <= (__read[155] ? __in : ((__apply_updates && __update_queue[155]) ? __l39_next[80][31:0] : __var[155]));
		__var[156][31:0] <= (__read[156] ? __in : ((__apply_updates && __update_queue[156]) ? __l39_next[81][31:0] : __var[156]));
		__var[157][31:0] <= (__read[157] ? __in : ((__apply_updates && __update_queue[157]) ? __l39_next[82][31:0] : __var[157]));
		__var[158][31:0] <= (__read[158] ? __in : ((__apply_updates && __update_queue[158]) ? __l39_next[83][31:0] : __var[158]));
		__var[159][31:0] <= (__read[159] ? __in : ((__apply_updates && __update_queue[159]) ? __l39_next[84][31:0] : __var[159]));
		__var[160][31:0] <= (__read[160] ? __in : ((__apply_updates && __update_queue[160]) ? __l39_next[85][31:0] : __var[160]));
		__var[161][31:0] <= (__read[161] ? __in : ((__apply_updates && __update_queue[161]) ? __l39_next[86][31:0] : __var[161]));
		__var[162][31:0] <= (__read[162] ? __in : ((__apply_updates && __update_queue[162]) ? __l39_next[87][31:0] : __var[162]));
		__var[163][31:0] <= (__read[163] ? __in : ((__apply_updates && __update_queue[163]) ? __l39_next[88][31:0] : __var[163]));
		__var[164][31:0] <= (__read[164] ? __in : ((__apply_updates && __update_queue[164]) ? __l39_next[89][31:0] : __var[164]));
		__var[165][31:0] <= (__read[165] ? __in : ((__apply_updates && __update_queue[165]) ? __l39_next[90][31:0] : __var[165]));
		__var[166][31:0] <= (__read[166] ? __in : ((__apply_updates && __update_queue[166]) ? __l39_next[91][31:0] : __var[166]));
		__var[167][31:0] <= (__read[167] ? __in : ((__apply_updates && __update_queue[167]) ? __l39_next[92][31:0] : __var[167]));
		__var[168][31:0] <= (__read[168] ? __in : ((__apply_updates && __update_queue[168]) ? __l39_next[93][31:0] : __var[168]));
		__var[169][31:0] <= (__read[169] ? __in : ((__apply_updates && __update_queue[169]) ? __l39_next[94][31:0] : __var[169]));
		__var[170][31:0] <= (__read[170] ? __in : ((__apply_updates && __update_queue[170]) ? __l39_next[95][31:0] : __var[170]));
		__var[171][31:0] <= (__read[171] ? __in : ((__apply_updates && __update_queue[171]) ? __l39_next[96][31:0] : __var[171]));
		__var[172][31:0] <= (__read[172] ? __in : ((__apply_updates && __update_queue[172]) ? __l39_next[97][31:0] : __var[172]));
		__var[173][31:0] <= (__read[173] ? __in : ((__apply_updates && __update_queue[173]) ? __l39_next[98][31:0] : __var[173]));
		__var[174][31:0] <= (__read[174] ? __in : ((__apply_updates && __update_queue[174]) ? __l39_next[99][31:0] : __var[174]));
		__var[175][31:0] <= (__read[175] ? __in : ((__apply_updates && __update_queue[175]) ? __l39_next[100][31:0] : __var[175]));
		__var[176][31:0] <= (__read[176] ? __in : ((__apply_updates && __update_queue[176]) ? __l39_next[101][31:0] : __var[176]));
		__var[177][31:0] <= (__read[177] ? __in : ((__apply_updates && __update_queue[177]) ? __l39_next[102][31:0] : __var[177]));
		__var[178][31:0] <= (__read[178] ? __in : ((__apply_updates && __update_queue[178]) ? __l39_next[103][31:0] : __var[178]));
		__var[179][31:0] <= (__read[179] ? __in : ((__apply_updates && __update_queue[179]) ? __l39_next[104][31:0] : __var[179]));
		__var[180][31:0] <= (__read[180] ? __in : ((__apply_updates && __update_queue[180]) ? __l39_next[105][31:0] : __var[180]));
		__var[181][31:0] <= (__read[181] ? __in : ((__apply_updates && __update_queue[181]) ? __l39_next[106][31:0] : __var[181]));
		__var[182][31:0] <= (__read[182] ? __in : ((__apply_updates && __update_queue[182]) ? __l39_next[107][31:0] : __var[182]));
		__var[183][31:0] <= (__read[183] ? __in : ((__apply_updates && __update_queue[183]) ? __l39_next[108][31:0] : __var[183]));
		__var[184][31:0] <= (__read[184] ? __in : ((__apply_updates && __update_queue[184]) ? __l39_next[109][31:0] : __var[184]));
		__var[185][31:0] <= (__read[185] ? __in : ((__apply_updates && __update_queue[185]) ? __l39_next[110][31:0] : __var[185]));
		__var[186][31:0] <= (__read[186] ? __in : ((__apply_updates && __update_queue[186]) ? __l39_next[111][31:0] : __var[186]));
		__var[187][31:0] <= (__read[187] ? __in : ((__apply_updates && __update_queue[187]) ? __l39_next[112][31:0] : __var[187]));
		__var[188][31:0] <= (__read[188] ? __in : ((__apply_updates && __update_queue[188]) ? __l39_next[113][31:0] : __var[188]));
		__var[189][31:0] <= (__read[189] ? __in : ((__apply_updates && __update_queue[189]) ? __l39_next[114][31:0] : __var[189]));
		__var[190][31:0] <= (__read[190] ? __in : ((__apply_updates && __update_queue[190]) ? __l39_next[115][31:0] : __var[190]));
		__var[191][31:0] <= (__read[191] ? __in : ((__apply_updates && __update_queue[191]) ? __l39_next[116][31:0] : __var[191]));
		__var[192][31:0] <= (__read[192] ? __in : ((__apply_updates && __update_queue[192]) ? __l39_next[117][31:0] : __var[192]));
		__var[193][31:0] <= (__read[193] ? __in : ((__apply_updates && __update_queue[193]) ? __l39_next[118][31:0] : __var[193]));
		__var[194][31:0] <= (__read[194] ? __in : ((__apply_updates && __update_queue[194]) ? __l39_next[119][31:0] : __var[194]));
		__var[195][31:0] <= (__read[195] ? __in : ((__apply_updates && __update_queue[195]) ? __l39_next[120][31:0] : __var[195]));
		__var[196][31:0] <= (__read[196] ? __in : ((__apply_updates && __update_queue[196]) ? __l39_next[121][31:0] : __var[196]));
		__var[197][31:0] <= (__read[197] ? __in : ((__apply_updates && __update_queue[197]) ? __l39_next[122][31:0] : __var[197]));
		__var[198][31:0] <= (__read[198] ? __in : ((__apply_updates && __update_queue[198]) ? __l39_next[123][31:0] : __var[198]));
		__var[199][31:0] <= (__read[199] ? __in : ((__apply_updates && __update_queue[199]) ? __l39_next[124][31:0] : __var[199]));
		__var[200][31:0] <= (__read[200] ? __in : ((__apply_updates && __update_queue[200]) ? __l39_next[125][31:0] : __var[200]));
		__var[201][31:0] <= (__read[201] ? __in : ((__apply_updates && __update_queue[201]) ? __l39_next[126][31:0] : __var[201]));
		__var[202][31:0] <= (__read[202] ? __in : ((__apply_updates && __update_queue[202]) ? __l39_next[127][31:0] : __var[202]));
		__var[203][31:0] <= (__read[203] ? __in : ((__apply_updates && __update_queue[203]) ? __l54_next[31:0] : __var[203]));
		__var[204][31:0] <= (__read[204] ? __in : ((__apply_updates && __update_queue[204]) ? __l64_next[0][31:0] : __var[204]));
		__var[205][31:0] <= (__read[205] ? __in : ((__apply_updates && __update_queue[205]) ? __l64_next[1][31:0] : __var[205]));
		__var[206][31:0] <= (__read[206] ? __in : ((__apply_updates && __update_queue[206]) ? __l64_next[2][31:0] : __var[206]));
		__var[207][31:0] <= (__read[207] ? __in : ((__apply_updates && __update_queue[207]) ? __l64_next[3][31:0] : __var[207]));
		__var[208][31:0] <= (__read[208] ? __in : ((__apply_updates && __update_queue[208]) ? __l64_next[4][31:0] : __var[208]));
		__var[209][31:0] <= (__read[209] ? __in : ((__apply_updates && __update_queue[209]) ? __l64_next[5][31:0] : __var[209]));
		__var[210][31:0] <= (__read[210] ? __in : ((__apply_updates && __update_queue[210]) ? __l64_next[6][31:0] : __var[210]));
		__var[211][31:0] <= (__read[211] ? __in : ((__apply_updates && __update_queue[211]) ? __l64_next[7][31:0] : __var[211]));
		__var[212][31:0] <= (__read[212] ? __in : ((__apply_updates && __update_queue[212]) ? __l64_next[8][31:0] : __var[212]));
		__var[213][31:0] <= (__read[213] ? __in : ((__apply_updates && __update_queue[213]) ? __l64_next[9][31:0] : __var[213]));
		__var[214][31:0] <= (__read[214] ? __in : ((__apply_updates && __update_queue[214]) ? __l64_next[10][31:0] : __var[214]));
		__var[215][31:0] <= (__read[215] ? __in : ((__apply_updates && __update_queue[215]) ? __l64_next[11][31:0] : __var[215]));
		__var[216][31:0] <= (__read[216] ? __in : ((__apply_updates && __update_queue[216]) ? __l64_next[12][31:0] : __var[216]));
		__var[217][31:0] <= (__read[217] ? __in : ((__apply_updates && __update_queue[217]) ? __l64_next[13][31:0] : __var[217]));
		__var[218][31:0] <= (__read[218] ? __in : ((__apply_updates && __update_queue[218]) ? __l64_next[14][31:0] : __var[218]));
		__var[219][31:0] <= (__read[219] ? __in : ((__apply_updates && __update_queue[219]) ? __l64_next[15][31:0] : __var[219]));
		__var[220][31:0] <= (__read[220] ? __in : ((__apply_updates && __update_queue[220]) ? __l64_next[16][31:0] : __var[220]));
		__var[221][31:0] <= (__read[221] ? __in : ((__apply_updates && __update_queue[221]) ? __l64_next[17][31:0] : __var[221]));
		__var[222][31:0] <= (__read[222] ? __in : ((__apply_updates && __update_queue[222]) ? __l64_next[18][31:0] : __var[222]));
		__var[223][31:0] <= (__read[223] ? __in : ((__apply_updates && __update_queue[223]) ? __l64_next[19][31:0] : __var[223]));
		__var[224][31:0] <= (__read[224] ? __in : ((__apply_updates && __update_queue[224]) ? __l64_next[20][31:0] : __var[224]));
		__var[225][31:0] <= (__read[225] ? __in : ((__apply_updates && __update_queue[225]) ? __l64_next[21][31:0] : __var[225]));
		__var[226][31:0] <= (__read[226] ? __in : ((__apply_updates && __update_queue[226]) ? __l64_next[22][31:0] : __var[226]));
		__var[227][31:0] <= (__read[227] ? __in : ((__apply_updates && __update_queue[227]) ? __l64_next[23][31:0] : __var[227]));
		__var[228][31:0] <= (__read[228] ? __in : ((__apply_updates && __update_queue[228]) ? __l64_next[24][31:0] : __var[228]));
		__var[229][31:0] <= (__read[229] ? __in : ((__apply_updates && __update_queue[229]) ? __l64_next[25][31:0] : __var[229]));
		__var[230][31:0] <= (__read[230] ? __in : ((__apply_updates && __update_queue[230]) ? __l64_next[26][31:0] : __var[230]));
		__var[231][31:0] <= (__read[231] ? __in : ((__apply_updates && __update_queue[231]) ? __l64_next[27][31:0] : __var[231]));
		__var[232][31:0] <= (__read[232] ? __in : ((__apply_updates && __update_queue[232]) ? __l64_next[28][31:0] : __var[232]));
		__var[233][31:0] <= (__read[233] ? __in : ((__apply_updates && __update_queue[233]) ? __l64_next[29][31:0] : __var[233]));
		__var[234][31:0] <= (__read[234] ? __in : ((__apply_updates && __update_queue[234]) ? __l64_next[30][31:0] : __var[234]));
		__var[235][31:0] <= (__read[235] ? __in : ((__apply_updates && __update_queue[235]) ? __l64_next[31][31:0] : __var[235]));
		__var[236][31:0] <= (__read[236] ? __in : ((__apply_updates && __update_queue[236]) ? __l75_next[31:0] : __var[236]));
		__var[237][31:0] <= (__read[237] ? __in : ((__apply_updates && __update_queue[237]) ? __l76_next[31:0] : __var[237]));
		if ((__apply_updates || __reset)) 
			__update_queue <= 0;
	end 
	always @(posedge __clk) begin
		if (__read[6]) 
			__feof[__in[6:1]] <= __in[0];
	end 
	reg[63:0] __out_buf_next[1:0];
	reg[63:0] __out_next;
	always @(posedge __clk) begin : __out_buf_block
		reg signed[31:0] t0;
		reg signed[31:0] t1;
		reg signed[31:0] t2;
		for (t0 = 0; (t0 <= 1); t0 = (t0 + 1)) begin
			__out_buf_next[t0] = 0;
		end 
		__out_buf_next[0] = (__out_buf_next[0] | (__write[0] ? __there_are_updates : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[2] ? __task_id[0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[5] ? __open_loop : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[7] ? __wait : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[8] ? __state[0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[9] ? __var[9][0:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[10] ? __var[10][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[11] ? __var[11][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[12] ? __var[12][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[13] ? __var[13][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[14] ? __var[14][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[15] ? __var[15][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[16] ? __var[16][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[17] ? __var[17][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[18] ? __var[18][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[19] ? __var[19][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[20] ? __var[20][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[21] ? __var[21][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[22] ? __var[22][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[23] ? __var[23][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[24] ? __var[24][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[25] ? __var[25][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[26] ? __var[26][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[27] ? __var[27][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[28] ? __var[28][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[29] ? __var[29][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[30] ? __var[30][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[31] ? __var[31][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[32] ? __var[32][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[33] ? __var[33][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[34] ? __var[34][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[35] ? __var[35][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[36] ? __var[36][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[37] ? __var[37][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[38] ? __var[38][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[39] ? __var[39][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[40] ? __var[40][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[41] ? __var[41][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[42] ? __var[42][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[43] ? __var[43][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[44] ? __var[44][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[45] ? __var[45][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[46] ? __var[46][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[47] ? __var[47][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[48] ? __var[48][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[49] ? __var[49][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[50] ? __var[50][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[51] ? __var[51][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[52] ? __var[52][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[53] ? __var[53][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[54] ? __var[54][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[55] ? __var[55][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[56] ? __var[56][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[57] ? __var[57][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[58] ? __var[58][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[59] ? __var[59][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[60] ? __var[60][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[61] ? __var[61][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[62] ? __var[62][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[63] ? __var[63][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[64] ? __var[64][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[65] ? __var[65][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[66] ? __var[66][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[67] ? __var[67][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[68] ? __var[68][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[69] ? __var[69][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[70] ? __var[70][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[71] ? __var[71][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[72] ? __var[72][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[73] ? __var[73][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[74] ? __var[74][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[75] ? __var[75][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[76] ? __var[76][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[77] ? __var[77][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[78] ? __var[78][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[79] ? __var[79][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[80] ? __var[80][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[81] ? __var[81][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[82] ? __var[82][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[83] ? __var[83][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[84] ? __var[84][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[85] ? __var[85][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[86] ? __var[86][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[87] ? __var[87][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[88] ? __var[88][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[89] ? __var[89][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[90] ? __var[90][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[91] ? __var[91][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[92] ? __var[92][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[93] ? __var[93][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[94] ? __var[94][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[95] ? __var[95][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[96] ? __var[96][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[97] ? __var[97][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[98] ? __var[98][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[99] ? __var[99][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[100] ? __var[100][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[101] ? __var[101][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[102] ? __var[102][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[103] ? __var[103][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[104] ? __var[104][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[105] ? __var[105][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[106] ? __var[106][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[107] ? __var[107][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[108] ? __var[108][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[109] ? __var[109][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[110] ? __var[110][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[111] ? __var[111][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[112] ? __var[112][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[113] ? __var[113][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[114] ? __var[114][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[115] ? __var[115][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[116] ? __var[116][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[117] ? __var[117][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[118] ? __var[118][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[119] ? __var[119][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[120] ? __var[120][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[121] ? __var[121][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[122] ? __var[122][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[123] ? __var[123][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[124] ? __var[124][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[125] ? __var[125][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[126] ? __var[126][31:0] : 0));
		__out_buf_next[0] = (__out_buf_next[0] | (__write[127] ? __var[127][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[128] ? __var[128][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[129] ? __var[129][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[130] ? __var[130][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[131] ? __var[131][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[132] ? __var[132][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[133] ? __var[133][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[134] ? __var[134][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[135] ? __var[135][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[136] ? __var[136][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[137] ? __var[137][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[138] ? __var[138][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[139] ? __var[139][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[140] ? __var[140][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[141] ? __var[141][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[142] ? __var[142][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[143] ? __var[143][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[144] ? __var[144][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[145] ? __var[145][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[146] ? __var[146][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[147] ? __var[147][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[148] ? __var[148][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[149] ? __var[149][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[150] ? __var[150][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[151] ? __var[151][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[152] ? __var[152][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[153] ? __var[153][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[154] ? __var[154][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[155] ? __var[155][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[156] ? __var[156][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[157] ? __var[157][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[158] ? __var[158][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[159] ? __var[159][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[160] ? __var[160][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[161] ? __var[161][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[162] ? __var[162][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[163] ? __var[163][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[164] ? __var[164][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[165] ? __var[165][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[166] ? __var[166][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[167] ? __var[167][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[168] ? __var[168][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[169] ? __var[169][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[170] ? __var[170][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[171] ? __var[171][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[172] ? __var[172][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[173] ? __var[173][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[174] ? __var[174][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[175] ? __var[175][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[176] ? __var[176][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[177] ? __var[177][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[178] ? __var[178][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[179] ? __var[179][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[180] ? __var[180][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[181] ? __var[181][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[182] ? __var[182][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[183] ? __var[183][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[184] ? __var[184][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[185] ? __var[185][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[186] ? __var[186][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[187] ? __var[187][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[188] ? __var[188][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[189] ? __var[189][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[190] ? __var[190][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[191] ? __var[191][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[192] ? __var[192][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[193] ? __var[193][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[194] ? __var[194][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[195] ? __var[195][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[196] ? __var[196][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[197] ? __var[197][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[198] ? __var[198][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[199] ? __var[199][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[200] ? __var[200][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[201] ? __var[201][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[202] ? __var[202][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[203] ? __var[203][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[204] ? __var[204][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[205] ? __var[205][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[206] ? __var[206][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[207] ? __var[207][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[208] ? __var[208][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[209] ? __var[209][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[210] ? __var[210][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[211] ? __var[211][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[212] ? __var[212][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[213] ? __var[213][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[214] ? __var[214][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[215] ? __var[215][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[216] ? __var[216][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[217] ? __var[217][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[218] ? __var[218][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[219] ? __var[219][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[220] ? __var[220][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[221] ? __var[221][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[222] ? __var[222][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[223] ? __var[223][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[224] ? __var[224][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[225] ? __var[225][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[226] ? __var[226][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[227] ? __var[227][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[228] ? __var[228][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[229] ? __var[229][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[230] ? __var[230][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[231] ? __var[231][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[232] ? __var[232][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[233] ? __var[233][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[234] ? __var[234][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[235] ? __var[235][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[236] ? __var[236][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[237] ? __var[237][31:0] : 0));
		__out_buf_next[1] = (__out_buf_next[1] | (__write[238] ? __l67[31:0] : 0));
		__out_next = 0;
		for (t2 = 0; (t2 <= 1); t2 = (t2 + 1)) begin
			__out_next = (__out_next | __out_buf[t2]);
		end 
		for (t1 = 0; (t1 <= 1); t1 = (t1 + 1)) begin
			__out_buf[t1] <= __out_buf_next[t1];
		end 
		__out <= __out_next;
		__out_valid_buf[3] <= (__in_valid & (!__in_read));
		__out_valid_buf[2] <= __out_valid_buf[3];
		__out_valid_buf[1] <= __out_valid_buf[2];
		__out_valid_buf[0] <= __out_valid_buf[1];
	end 
	assign __out_data = __out;
	assign __out_valid = __out_valid_buf[0];
	assign __wait = ((__open_loop_tick || __any_triggers) || ((!__all_final) && (!__there_were_tasks)));
endmodule

module program_logic(
  input wire clk,
  input wire reset,

  input wire         softreg_req_valid,
  input wire         softreg_req_isWrite,
  input wire[31:0]   softreg_req_addr,
  input wire[63:0]   softreg_req_data,

  output wire        softreg_resp_valid,
  output wire[63:0]  softreg_resp_data
);

  parameter app_num = 0;

  // Register module signals
  reg        valid_in;
  reg        write_in;
  reg        read_in;
  reg[13:0]  addr_in;
  reg[63:0]  data_in;

  wire       valid_out;
  wire[63:0] data_out;
  reg        valid_out_reg;
  reg[63:0]  data_out_reg;

  always @(posedge clk) begin
    if (reset) begin
      valid_in <= 1'b0;
      write_in <= 1'b0;
      read_in <= 1'b0;
      addr_in <= 14'b0;
      data_in <= 64'b0;
    end else begin
      valid_in <= softreg_req_valid;
      write_in <= softreg_req_valid & softreg_req_isWrite;
      read_in <= softreg_req_valid & ~softreg_req_isWrite;
      addr_in <= softreg_req_addr[16:3];
      data_in <= softreg_req_data;
    end

    if (reset) begin
      valid_out_reg <= 1'b0;
      data_out_reg <= 64'b0;
    end else begin
      valid_out_reg <= valid_out;
      data_out_reg <= data_out;
    end
  end

  assign softreg_resp_valid = valid_out_reg;
  assign softreg_resp_data = data_out_reg;

  // Module Instantiations:
  generate
  if (app_num == 0) begin
    M0 m (
      .__clk(clk),
      .__in_read(write_in),
      .__in_vid(addr_in),
      .__in_data(data_in),
      .__in_valid(valid_in),
      .__out_data(data_out),
      .__out_valid(valid_out)
    );
  end
  endgenerate
endmodule
